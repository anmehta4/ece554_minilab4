module memA
#(
  parameter BITS_AB=8,
  parameter DIM=8
)
(
  input clk,rst_n,en,WrEn,
  input signed [BITS_AB-1:0] Ain [DIM-1:0],
  input [$clog2(DIM)-1:0] Arow,
  output signed [BITS_AB-1:0] Aout [DIM-1:0]
);



endmodule
